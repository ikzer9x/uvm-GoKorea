   //---------------------------------------------------------------------------
   // Typedef: coasia_sequencer
   //--------------------------------------------------------------------------- 
   typedef uvm_sequencer#(coasia_transaction) coasia_sequencer; 
